`timescale 1ns / 1ps
/*
 * Copyright (c) 2023 Govardhan
 *
 * Permission is hereby granted, free of charge, to any person obtaining a copy
 * of this software and associated documentation files (the "Software"), to deal
 * in the Software without restriction, including without limitation the rights
 * to use, copy, modify, merge, publish, distribute, sublicense, and/or sell
 * copies of the Software, and to permit persons to whom the Software is
 * furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included in
 * all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS OR
 * IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL THE
 * AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM,
 * OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN
 * THE SOFTWARE.
 */

module Single_Cycle_Core(
    input  wire        clk, reset,
    input  wire [31:0] Instr,
    input  wire [31:0] ReadData,
    output wire [31:0] PC,
    output wire        MemWrite,
    output wire [31:0] ALUResult,
    output wire [31:0] WriteData
);

    wire        ALUSrc, RegWrite, Jump, Branch;
    wire        PCSrc; // not used at top-level now, kept for compatibility
    wire [1:0]  ResultSrc, ImmSrc;
    wire [3:0]  ALUControl;
	wire MemRead;

    // instantiate control unit (export Branch, Jump to datapath)
    Control_Unit Control (
        .op(Instr[6:0]),
        .funct3(Instr[14:12]),
        .funct7b5(Instr[30]),
        .Zero(),               // datapath drives Zero, keep wire unused here
        .ResultSrc(ResultSrc),
        .MemWrite(MemWrite),
		.MemRead(MemRead),
        .PCSrc(PCSrc),
        .ALUSrc(ALUSrc),
        .RegWrite(RegWrite),
        .Branch(Branch),
        .Jump(Jump),
        .ImmSrc(ImmSrc),
        .ALUControl(ALUControl)
    );

    // Instantiate the datapath with named port mapping to avoid positional mismatch
    Core_Datapath Datapath (
        .clk(clk),
        .reset(reset),
        .ResultSrc(ResultSrc),
        .PCSrc(PCSrc),         // still present in datapath ports (unused internally)
        .ALUSrc(ALUSrc),
        .RegWrite(RegWrite),
        .ImmSrc(ImmSrc),
        .ALUControl(ALUControl),
        .Instr(Instr),         // IF-stage Instr from IMEM
        .ReadData(ReadData),
        .Branch(Branch),
        .Jump(Jump),
		.MemWrite(MemWrite),
		.MemRead(MemRead),
        .Zero(),               // datapath outputs Zero internally; not used at top-level
        .PC(PC),
        .ALUResult(ALUResult),
        .WriteData(WriteData)
    );

endmodule
